module test ();

  initial begin

    $display("Hello");

  end

  string name = "Aizaz";
  
  initial begin
    $display(name);
  end
endmodule
