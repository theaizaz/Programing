module test ();

  initial begin

    $display("Hello");

  end

	string fname = "Aizaz";
  	string lname = "khan";
  
  initial begin
    
    $display("Hello %s ",fname);
    
  end
endmodule
